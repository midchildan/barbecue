// barbecue - a simple processor based on RISC-V
// Copyright © 2017 Team Barbecue
//
// Permission is hereby granted, free of charge, to any person obtaining
// a copy of this software and associated documentation files (the "Software"),
// to deal in the Software without restriction, including without limitation
// the rights to use, copy, modify, merge, publish, distribute, sublicense,
// and/or sell copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included
// in all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
// OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM,
// DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
// TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE
// OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.


module top (
  input clk,
  input reset
);

  `include "constants.vh"

  wire [XLEN-1:0] imem_addr;
  wire [XLEN-1:0] imem_rdata;
  wire [XLEN-1:0] dmem_addr;
  wire [XLEN-1:0] dmem_rdata;
  wire [XLEN-1:0] dmem_wdata;
  wire dmem_we;

  datapath datapath (
    // input
    .clk(clk),
    .reset(reset),
    .imem_rdata(imem_rdata),
    .dmem_rdata(dmem_rdata),

    // output
    .imem_addr(imem_addr),
    .dmem_addr(dmem_addr),
    .dmem_wdata(dmem_wdata),
    .dmem_we(dmem_we)
  );

  imem imem (
    // input
    .clk(clk),
    .addr(imem_addr),

    // output
    .rdata(imem_rdata)
  );

  dmem dmem (
    // input
    .clk(clk),
    .addr(dmem_addr),
    .wdata(dmem_wdata),
    .we(dmem_we),

    // output
    .rdata(dmem_rdata)
  );

endmodule
